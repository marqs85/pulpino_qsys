`ifndef ADBG_CONFIG_SV
`define ADBG_CONFIG_SV

//`define ENABLE_ADV_DBG_IF
//`define DBG_WISHBONE_SUPPORTED

`endif
